`ifndef ADDER_SEQUENCER_SV
`define ADDER_SEQUENCER_SV

typedef uvm_sequencer #(adder_sequence_item) adder_sequencer;

`endif // ADDER_SEQUENCER_SV
