`ifndef TOP_TEST_PKG_SV
`define TOP_TEST_PKG_SV

package top_test_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "top_test.sv"

endpackage : top_test_pkg

`endif // TOP_TEST_PKG_SV
