`ifndef ADDER_TYPEDEFS_SV
`define ADDER_TYPEDEFS_SV

typedef enum {TRANS_FISRT, TRANS_MIDDLE, TRANS_LAST} trans_stage_t;
typedef enum {TRANS_SYNC,  TRANS_ASYNC} trans_type_t;

`endif // ADDER_TYPEDEFS_SV
